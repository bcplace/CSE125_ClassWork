module palindrome
  #(parameter [31:0] depth_p = 32'd10)
   (input [0:0] clk_i
   ,input [0:0] reset_i
   ,input [3:0] symbol_i
   ,input [0:0] valid_i
   ,output [0:0] overflow_o // Not required, but provided for debugging
   ,output [0:0] palindrome_o);

   // Your code here:
     
       
endmodule


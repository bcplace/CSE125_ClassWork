module multiplier
  #(parameter width_p = 8)
  (input [width_p - 1:0]  a_i,
   input [width_p - 1:0]  b_i, 
   output [(2*width_p) - 1:0] prod_o);

   assign prod_o = (a_i * b_i);

   // Write your immediate and concurrent assertions here

   // The synthesized code below does not implement the correct
   // behavior (but the error is simple).
   // 
   // You must write two concurrent assertions, one demonstrating your understanding
   //
   //  - One must fail (Demonstrating your understanding of how to
   //  write a concurrent assertion that checks for correct behavior.)
   //
   //  - One must pass (Demonstrating your understanding of the bug)
   //

   // Use `ifdef FORMAL to hide your concurrent assertion from iverilog
`ifdef FORMAL

`endif

endmodule

module multiplier_synth
  #(parameter width_p = 8)
  (input [width_p - 1:0]  a_i,
   input [width_p - 1:0]  b_i, 
   output [(2*width_p) - 1:0] prod_o);

   // Write your immediate and concurrent assertions here
   
   // The synthesized code below does not implement the correct
   // behavior (but the error is simple).
   // 
   // You must write two concurrent assertions, one demonstrating your understanding
   //
   //  - One must fail (Demonstrating your understanding of how to
   //  write a concurrent assertion that checks for correct behavior.)
   //
   //  - One must pass (Demonstrating your understanding of the bug)
   //

   // Use `ifdef FORMAL to hide your concurrent assertion from iverilog
`ifdef FORMAL

`endif

   yosys_multiplier
     #()
   mul_synth_i
     (.a_i(a_i)
     ,.b_i(b_i)
     ,.prod_o(prod_o));

endmodule

(* hdlname = "\\multiplier" *)
(* dynports =  1  *)
(* top =  1  *)
(* src = "multiplier.sv:1.1-9.10" *)
module yosys_multiplier(a_i, b_i, prod_o);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  wire _192_;
  wire _193_;
  wire _194_;
  wire _195_;
  wire _196_;
  wire _197_;
  wire _198_;
  wire _199_;
  wire _200_;
  wire _201_;
  wire _202_;
  wire _203_;
  wire _204_;
  wire _205_;
  wire _206_;
  wire _207_;
  wire _208_;
  wire _209_;
  wire _210_;
  wire _211_;
  wire _212_;
  wire _213_;
  wire _214_;
  wire _215_;
  wire _216_;
  wire _217_;
  wire _218_;
  wire _219_;
  wire _220_;
  wire _221_;
  wire _222_;
  wire _223_;
  wire _224_;
  wire _225_;
  wire _226_;
  wire _227_;
  wire _228_;
  wire _229_;
  wire _230_;
  wire _231_;
  wire _232_;
  wire _233_;
  wire _234_;
  wire _235_;
  wire _236_;
  wire _237_;
  wire _238_;
  wire _239_;
  wire _240_;
  wire _241_;
  wire _242_;
  wire _243_;
  wire _244_;
  wire _245_;
  wire _246_;
  wire _247_;
  wire _248_;
  wire _249_;
  wire _250_;
  wire _251_;
  wire _252_;
  wire _253_;
  wire _254_;
  wire _255_;
  wire _256_;
  wire _257_;
  wire _258_;
  wire _259_;
  wire _260_;
  wire _261_;
  wire _262_;
  wire _263_;
  wire _264_;
  wire _265_;
  wire _266_;
  wire _267_;
  wire _268_;
  wire _269_;
  wire _270_;
  wire _271_;
  wire _272_;
  wire _273_;
  wire _274_;
  wire _275_;
  wire _276_;
  wire _277_;
  wire _278_;
  wire _279_;
  wire _280_;
  wire _281_;
  wire _282_;
  wire _283_;
  wire _284_;
  wire _285_;
  wire _286_;
  wire _287_;
  wire _288_;
  wire _289_;
  wire _290_;
  wire _291_;
  wire _292_;
  wire _293_;
  wire _294_;
  wire _295_;
  wire _296_;
  wire _297_;
  wire _298_;
  wire _299_;
  wire _300_;
  wire _301_;
  wire _302_;
  wire _303_;
  wire _304_;
  wire _305_;
  wire _306_;
  wire _307_;
  wire _308_;
  wire _309_;
  wire _310_;
  wire _311_;
  wire _312_;
  wire _313_;
  wire _314_;
  wire _315_;
  wire _316_;
  wire _317_;
  wire _318_;
  wire _319_;
  wire _320_;
  wire _321_;
  wire _322_;
  wire _323_;
  wire _324_;
  wire _325_;
  wire _326_;
  wire _327_;
  wire _328_;
  wire _329_;
  wire _330_;
  wire _331_;
  wire _332_;
  wire _333_;
  wire _334_;
  (* src = "multiplier.sv:3.27-3.30" *)
  input [7:0] a_i;
  wire [7:0] a_i;
  (* src = "multiplier.sv:4.27-4.30" *)
  input [7:0] b_i;
  wire [7:0] b_i;
  (* src = "multiplier.sv:5.31-5.37" *)
  output [15:0] prod_o;
  wire [15:0] prod_o;
  assign _300_ = _283_ & ~(_284_);
  assign _301_ = _299_ & ~(_300_);
  assign _302_ = _301_ ^ _298_;
  assign _303_ = b_i[3] & a_i[1];
  assign _304_ = b_i[4] & a_i[0];
  assign _305_ = ~(_304_ ^ _303_);
  assign _306_ = _305_ ^ _302_;
  assign _307_ = _288_ | _285_;
  assign _308_ = _289_ & ~(_291_);
  assign _309_ = _307_ & ~(_308_);
  assign _310_ = ~(_309_ ^ _306_);
  assign _311_ = _293_ & ~(_292_);
  assign prod_o[4] = ~(_311_ ^ _310_);
  assign _312_ = ~(a_i[6] & b_i[0]);
  assign _313_ = ~(b_i[1] & a_i[5]);
  assign _314_ = _313_ ^ _312_;
  assign _315_ = ~(b_i[2] & a_i[4]);
  assign _316_ = _315_ ^ _314_;
  assign _317_ = ~(a_i[5] & b_i[0]);
  assign _318_ = b_i[1] & a_i[4];
  assign _319_ = _317_ | ~(_318_);
  assign _320_ = b_i[2] & a_i[3];
  assign _321_ = _318_ ^ _317_;
  assign _322_ = _320_ & ~(_321_);
  assign _323_ = _319_ & ~(_322_);
  assign _324_ = _323_ ^ _316_;
  assign _325_ = b_i[3] & a_i[3];
  assign _326_ = b_i[4] & a_i[2];
  assign _327_ = _326_ ^ _325_;
  assign _328_ = ~(b_i[5] & a_i[1]);
  assign _329_ = _328_ ^ _327_;
  assign _330_ = _329_ ^ _324_;
  assign _331_ = ~(_321_ ^ _320_);
  assign _332_ = _295_ | _294_;
  assign _333_ = _296_ & ~(_297_);
  assign _334_ = _332_ & ~(_333_);
  assign _000_ = _334_ | ~(_331_);
  assign _001_ = b_i[3] & a_i[2];
  assign _002_ = b_i[4] & a_i[1];
  assign _003_ = _002_ ^ _001_;
  assign _004_ = b_i[5] & a_i[0];
  assign _005_ = _004_ ^ _003_;
  assign _006_ = _334_ ^ _331_;
  assign _007_ = _005_ & ~(_006_);
  assign _008_ = _000_ & ~(_007_);
  assign _009_ = _008_ ^ _330_;
  assign _010_ = ~(_002_ & _001_);
  assign _011_ = _004_ & _003_;
  assign _012_ = _010_ & ~(_011_);
  assign _013_ = b_i[6] & a_i[0];
  assign _014_ = _013_ ^ _012_;
  assign _015_ = ~(_014_ ^ _009_);
  assign _016_ = ~(_006_ ^ _005_);
  assign _017_ = _301_ | _298_;
  assign _018_ = _302_ & ~(_305_);
  assign _019_ = _017_ & ~(_018_);
  assign _020_ = _019_ | ~(_016_);
  assign _021_ = _304_ & _303_;
  assign _022_ = _019_ ^ _016_;
  assign _023_ = _021_ & ~(_022_);
  assign _024_ = _020_ & ~(_023_);
  assign _025_ = _024_ ^ _015_;
  assign _026_ = _022_ ^ _021_;
  assign _027_ = _309_ | _306_;
  assign _028_ = _027_ | _026_;
  assign _029_ = ~(_028_ ^ _025_);
  assign _030_ = _027_ ^ _026_;
  assign _031_ = _311_ & ~(_310_);
  assign _032_ = _031_ & _030_;
  assign prod_o[6] = ~(_032_ ^ _029_);
  assign _033_ = ~(a_i[7] & b_i[0]);
  assign _034_ = ~(b_i[1] & a_i[6]);
  assign _035_ = _034_ ^ _033_;
  assign _036_ = ~(b_i[2] & a_i[5]);
  assign _037_ = _036_ ^ _035_;
  assign _038_ = _313_ | _312_;
  assign _039_ = _314_ & ~(_315_);
  assign _040_ = _038_ & ~(_039_);
  assign _041_ = _040_ ^ _037_;
  assign _042_ = b_i[3] & a_i[4];
  assign _043_ = b_i[4] & a_i[3];
  assign _044_ = _043_ ^ _042_;
  assign _045_ = ~(b_i[5] & a_i[2]);
  assign _046_ = _045_ ^ _044_;
  assign _047_ = _046_ ^ _041_;
  assign _048_ = _323_ | _316_;
  assign _049_ = _324_ & ~(_329_);
  assign _050_ = _048_ & ~(_049_);
  assign _051_ = _050_ ^ _047_;
  assign _052_ = ~(_326_ & _325_);
  assign _053_ = _327_ & ~(_328_);
  assign _054_ = _052_ & ~(_053_);
  assign _055_ = b_i[6] & a_i[1];
  assign _056_ = ~_055_;
  assign _057_ = _056_ ^ _054_;
  assign _058_ = b_i[7] & a_i[0];
  assign _059_ = ~_058_;
  assign _060_ = _059_ ^ _057_;
  assign _061_ = _060_ ^ _051_;
  assign _062_ = _008_ | _330_;
  assign _063_ = _009_ & ~(_014_);
  assign _064_ = _062_ & ~(_063_);
  assign _065_ = _064_ ^ _061_;
  assign _066_ = _013_ & ~(_012_);
  assign _067_ = ~_066_;
  assign _068_ = _067_ ^ _065_;
  assign _069_ = _015_ & ~(_024_);
  assign _070_ = _069_ ^ _068_;
  assign _071_ = _028_ | _025_;
  assign _072_ = _032_ & ~(_029_);
  assign _073_ = _071_ & ~(_072_);
  assign prod_o[7] = _073_ ^ _070_;
  assign _074_ = ~(b_i[1] & a_i[7]);
  assign _075_ = b_i[2] & a_i[6];
  assign _076_ = _075_ ^ _074_;
  assign _077_ = _034_ | _033_;
  assign _078_ = _035_ & ~(_036_);
  assign _079_ = _077_ & ~(_078_);
  assign _080_ = _079_ ^ _076_;
  assign _081_ = b_i[3] & a_i[5];
  assign _082_ = b_i[4] & a_i[4];
  assign _083_ = _082_ ^ _081_;
  assign _084_ = ~(b_i[5] & a_i[3]);
  assign _085_ = _084_ ^ _083_;
  assign _086_ = _085_ ^ _080_;
  assign _087_ = _040_ | _037_;
  assign _088_ = _041_ & ~(_046_);
  assign _089_ = _087_ & ~(_088_);
  assign _090_ = _089_ ^ _086_;
  assign _091_ = ~(_043_ & _042_);
  assign _092_ = _044_ & ~(_045_);
  assign _093_ = _091_ & ~(_092_);
  assign _094_ = b_i[6] & a_i[2];
  assign _095_ = _094_ ^ _093_;
  assign _096_ = b_i[7] & a_i[1];
  assign _097_ = _096_ ^ _095_;
  assign _098_ = _097_ ^ _090_;
  assign _099_ = _050_ | _047_;
  assign _100_ = _051_ & ~(_060_);
  assign _101_ = _099_ & ~(_100_);
  assign _102_ = _101_ ^ _098_;
  assign _103_ = _056_ | _054_;
  assign _104_ = _057_ & ~(_059_);
  assign _105_ = _103_ & ~(_104_);
  assign _106_ = _105_ ^ _102_;
  assign _107_ = _064_ | _061_;
  assign _108_ = _065_ & ~(_067_);
  assign _109_ = _107_ & ~(_108_);
  assign _110_ = ~(_109_ ^ _106_);
  assign _111_ = _068_ | ~(_069_);
  assign _112_ = ~(_071_ | _070_);
  assign _113_ = _111_ & ~(_112_);
  assign _114_ = _070_ | _029_;
  assign _115_ = _032_ & ~(_114_);
  assign _116_ = _113_ & ~(_115_);
  assign prod_o[8] = _116_ ^ _110_;
  assign _117_ = b_i[2] & a_i[7];
  assign _118_ = _075_ & ~(_074_);
  assign _119_ = _118_ ^ _117_;
  assign _120_ = b_i[3] & a_i[6];
  assign _121_ = b_i[4] & a_i[5];
  assign _122_ = _121_ ^ _120_;
  assign _123_ = b_i[5] & a_i[4];
  assign _124_ = ~_123_;
  assign _125_ = _124_ ^ _122_;
  assign _126_ = _125_ ^ _119_;
  assign _127_ = _079_ | _076_;
  assign _128_ = _080_ & ~(_085_);
  assign _129_ = _127_ & ~(_128_);
  assign _130_ = _129_ ^ _126_;
  assign _131_ = ~(_082_ & _081_);
  assign _132_ = _083_ & ~(_084_);
  assign _133_ = _131_ & ~(_132_);
  assign _134_ = b_i[6] & a_i[3];
  assign _135_ = _134_ ^ _133_;
  assign _136_ = b_i[7] & a_i[2];
  assign _137_ = _136_ ^ _135_;
  assign _138_ = _137_ ^ _130_;
  assign _139_ = _089_ | _086_;
  assign _140_ = _090_ & ~(_097_);
  assign _141_ = _139_ & ~(_140_);
  assign _142_ = _141_ ^ _138_;
  assign _143_ = _093_ | ~(_094_);
  assign _144_ = _096_ & ~(_095_);
  assign _145_ = _143_ & ~(_144_);
  assign _146_ = ~(_145_ ^ _142_);
  assign _147_ = _101_ | _098_;
  assign _148_ = _102_ & ~(_105_);
  assign _149_ = _147_ & ~(_148_);
  assign _150_ = _149_ ^ _146_;
  assign _151_ = _109_ | _106_;
  assign _152_ = _115_ | ~(_113_);
  assign _153_ = _152_ & ~(_110_);
  assign _154_ = _151_ & ~(_153_);
  assign prod_o[9] = _154_ ^ _150_;
  assign _155_ = b_i[3] & a_i[7];
  assign _156_ = b_i[4] & a_i[6];
  assign _157_ = ~(_156_ ^ _155_);
  assign _158_ = b_i[5] & a_i[5];
  assign _159_ = _158_ ^ _157_;
  assign _160_ = ~(_118_ & _117_);
  assign _161_ = _119_ & ~(_125_);
  assign _162_ = _160_ & ~(_161_);
  assign _163_ = _162_ ^ _159_;
  assign _164_ = _121_ & _120_;
  assign _165_ = _122_ & ~(_124_);
  assign _166_ = ~(_165_ | _164_);
  assign _167_ = b_i[6] & a_i[4];
  assign _168_ = _167_ ^ _166_;
  assign _169_ = b_i[7] & a_i[3];
  assign _170_ = _169_ ^ _168_;
  assign _171_ = _170_ ^ _163_;
  assign _172_ = _129_ | _126_;
  assign _173_ = _130_ & ~(_137_);
  assign _174_ = _172_ & ~(_173_);
  assign _175_ = _174_ ^ _171_;
  assign _176_ = _133_ | ~(_134_);
  assign _177_ = _136_ & ~(_135_);
  assign _178_ = _176_ & ~(_177_);
  assign _179_ = _178_ ^ _175_;
  assign _180_ = _141_ | _138_;
  assign _181_ = _142_ & ~(_145_);
  assign _182_ = _180_ & ~(_181_);
  assign _183_ = ~(_182_ ^ _179_);
  assign _184_ = _149_ | ~(_146_);
  assign _185_ = ~(_151_ | _150_);
  assign _186_ = _185_ | ~(_184_);
  assign _187_ = _150_ | _110_;
  assign _188_ = _187_ | _116_;
  assign _189_ = _188_ & ~(_186_);
  assign prod_o[10] = _189_ ^ _183_;
  assign _190_ = b_i[4] & a_i[7];
  assign _191_ = b_i[5] & a_i[6];
  assign _192_ = ~(_191_ ^ _190_);
  assign _193_ = ~_192_;
  assign _194_ = _156_ & _155_;
  assign _195_ = _158_ & ~(_157_);
  assign _196_ = ~(_195_ | _194_);
  assign _197_ = b_i[6] & a_i[5];
  assign _198_ = _197_ ^ _196_;
  assign _199_ = b_i[7] & a_i[4];
  assign _200_ = _199_ ^ _198_;
  assign _201_ = _200_ ^ _193_;
  assign _202_ = _162_ | _159_;
  assign _203_ = _163_ & ~(_170_);
  assign _204_ = _202_ & ~(_203_);
  assign _205_ = _204_ ^ _201_;
  assign _206_ = _166_ | ~(_167_);
  assign _207_ = _169_ & ~(_168_);
  assign _208_ = _206_ & ~(_207_);
  assign _209_ = _208_ ^ _205_;
  assign _210_ = _174_ | _171_;
  assign _211_ = _175_ & ~(_178_);
  assign _212_ = _210_ & ~(_211_);
  assign _213_ = ~(_212_ ^ _209_);
  assign _214_ = _182_ | _179_;
  assign _215_ = ~(_189_ | _183_);
  assign _216_ = _214_ & ~(_215_);
  assign prod_o[11] = _216_ ^ _213_;
  assign _217_ = b_i[5] & a_i[7];
  assign _218_ = _191_ & _190_;
  assign _219_ = b_i[6] & a_i[6];
  assign _220_ = ~(_219_ ^ _218_);
  assign _221_ = b_i[7] & a_i[5];
  assign _222_ = _221_ ^ _220_;
  assign _223_ = _222_ ^ _217_;
  assign _224_ = _193_ & ~(_200_);
  assign _225_ = _224_ ^ _223_;
  assign _226_ = _196_ | ~(_197_);
  assign _227_ = _199_ & ~(_198_);
  assign _228_ = _226_ & ~(_227_);
  assign _229_ = ~(_228_ ^ _225_);
  assign _230_ = _204_ | _201_;
  assign _231_ = _205_ & ~(_208_);
  assign _232_ = _230_ & ~(_231_);
  assign _233_ = ~(_232_ ^ _229_);
  assign _235_ = _212_ | _209_;
  assign _236_ = ~(_214_ | _213_);
  assign _237_ = _235_ & ~(_236_);
  assign _238_ = _213_ | _183_;
  assign _239_ = _186_ & ~(_238_);
  assign _240_ = _237_ & ~(_239_);
  assign _241_ = _238_ | _187_;
  assign _242_ = _152_ & ~(_241_);
  assign _243_ = _240_ & ~(_242_);
  assign prod_o[12] = _243_ ^ _233_;
  assign _245_ = b_i[6] & a_i[7];
  assign _246_ = b_i[7] & a_i[6];
  assign _247_ = ~(_246_ ^ _245_);
  assign _248_ = _217_ & ~(_222_);
  assign _249_ = _248_ ^ _247_;
  assign _250_ = ~(_219_ & _218_);
  assign _251_ = _221_ & ~(_220_);
  assign _252_ = _250_ & ~(_251_);
  assign _253_ = ~(_252_ ^ _249_);
  assign _254_ = _223_ | ~(_224_);
  assign _255_ = ~(_228_ | _225_);
  assign _256_ = _254_ & ~(_255_);
  assign _257_ = ~(_256_ ^ _253_);
  assign _258_ = _232_ | _229_;
  assign _259_ = ~(_243_ | _233_);
  assign _260_ = _258_ & ~(_259_);
  assign prod_o[13] = _260_ ^ _257_;
  assign _261_ = b_i[7] & a_i[7];
  assign _262_ = _246_ & _245_;
  assign _263_ = _262_ ^ _261_;
  assign _265_ = _247_ | ~(_248_);
  assign _266_ = ~(_252_ | _249_);
  assign _267_ = _265_ & ~(_266_);
  assign _268_ = _267_ ^ _263_;
  assign _269_ = _256_ | _253_;
  assign _270_ = ~(_258_ | _257_);
  assign _271_ = _269_ & ~(_270_);
  assign _272_ = _257_ | _233_;
  assign _273_ = ~(_272_ | _243_);
  assign _274_ = _271_ & ~(_273_);
  assign prod_o[14] = _274_ ^ _268_;
  assign prod_o[5] = _031_ ^ _030_;
  assign prod_o[0] = b_i[0] & a_i[0];
  assign _234_ = a_i[1] & b_i[0];
  assign _244_ = b_i[1] & a_i[0];
  assign prod_o[1] = _244_ ^ _234_;
  assign _264_ = a_i[2] & b_i[0];
  assign _275_ = b_i[1] & a_i[1];
  assign _276_ = _275_ ^ _264_;
  assign _277_ = b_i[2] & a_i[0];
  assign _278_ = ~_277_;
  assign _279_ = _278_ ^ _276_;
  assign _280_ = _244_ & _234_;
  assign prod_o[2] = ~(_280_ ^ _279_);
  assign _281_ = ~(a_i[3] & b_i[0]);
  assign _282_ = ~(b_i[1] & a_i[2]);
  assign _283_ = _282_ ^ _281_;
  assign _284_ = ~(b_i[2] & a_i[1]);
  assign _285_ = _284_ ^ _283_;
  assign _286_ = ~(_275_ & _264_);
  assign _287_ = _276_ & ~(_278_);
  assign _288_ = _286_ & ~(_287_);
  assign _289_ = _288_ ^ _285_;
  assign _290_ = b_i[3] & a_i[0];
  assign _291_ = ~_290_;
  assign _292_ = _291_ ^ _289_;
  assign _293_ = _280_ & ~(_279_);
  assign prod_o[3] = ~(_293_ ^ _292_);
  assign _294_ = ~(a_i[4] & b_i[0]);
  assign _295_ = ~(b_i[1] & a_i[3]);
  assign _296_ = _295_ ^ _294_;
  assign _297_ = ~(b_i[2] & a_i[2]);
  assign _298_ = _297_ ^ _296_;
  assign _299_ = _282_ | _281_;
  assign prod_o[15] = 1'h0;
endmodule

module countones
  #(parameter width_p = 32)
  (input [width_p - 1:0] binary_i
  ,output [$clog2(width_p) :0] count_o);

  logic [$clog2(width_p) :0] count_l; 

  // For extra credit (25% of Lab 3/Part 3): 
  // 
  // Re-write this loop to synthesize into better hardware. You may
  // not use the $countones() function (though it is synthesizable).
  // 
  // Demonstrate your improvement using the Yosys commands in Piazza.
  always_comb begin
     count_l = 0;
     for(logic [31:0] i = 0; i < width_p; i++) begin
        count_l += {{$clog2(width_p-1){1'b0}},binary_i[i]};
     end
  end
  assign count_o = count_l;

  // Write your immediate and concurrent assertions here

  // The synthesized code below does not implement the correct
  // behavior (but the error is simple).
  // 
  // You must write two concurrent assertions, one demonstrating your understanding
  //
  //  - One must fail (Demonstrating your understanding of how to
  //  write a concurrent assertion that checks for correct behavior.)
  //
  //  - One must pass (Demonstrating your understanding of the bug)
  //

  // Use `ifdef FORMAL to hide your concurrent assertion from iverilog
`ifdef FORMAL

`endif

endmodule

module countones_synth
  #(parameter width_p = 32)
  (input [width_p - 1:0] binary_i
  ,output [$clog2(width_p) :0] count_o);

  // Write your immediate and concurrent assertions here

  // The synthesized code below does not implement the correct
  // behavior (but the error is simple).
  // 
  // You must write two concurrent assertions, one demonstrating your understanding
  //
  //  - One must fail (Demonstrating your understanding of how to
  //  write a concurrent assertion that checks for correct behavior.)
  //
  //  - One must pass (Demonstrating your understanding of the bug)
  //

  // Use `ifdef FORMAL to hide your concurrent assertion from iverilog
`ifdef FORMAL

`endif

  yosys_countones
    #()
  countones_synth_i
    (.binary_i(binary_i)
    ,.count_o(count_o));

endmodule


/* Generated by Yosys 0.25 (git sha1 e02b7f64bc7, clang 14.0.0 -fPIC -Os) */

(* hdlname = "\\countones" *)
(* dynports =  1  *)
(* top =  1  *)
(* src = "countones.sv:1.1-43.10" *)
module yosys_countones(binary_i, count_o);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  (* src = "countones.sv:3.26-3.34" *)
  input [31:0] binary_i;
  wire [31:0] binary_i;
  (* src = "countones.sv:4.32-4.39" *)
  output [5:0] count_o;
  wire [5:0] count_o;
  assign _133_ = _126_ ^ _125_;
  assign _134_ = ~(_133_ ^ binary_i[2]);
  assign _135_ = _134_ ^ binary_i[1];
  assign _136_ = ~(_131_ ^ binary_i[12]);
  assign _137_ = _135_ & ~(_136_);
  assign _138_ = _132_ & ~(_137_);
  assign _139_ = _138_ ^ _130_;
  assign _140_ = _133_ | binary_i[2];
  assign _141_ = ~(_134_ | binary_i[1]);
  assign _000_ = _140_ & ~(_141_);
  assign _001_ = binary_i[6] | binary_i[5];
  assign _002_ = ~(_124_ | binary_i[7]);
  assign _003_ = _001_ & ~(_002_);
  assign _004_ = _003_ ^ _000_;
  assign _005_ = binary_i[15] | binary_i[11];
  assign _006_ = ~binary_i[8];
  assign _007_ = ~(binary_i[15] ^ binary_i[11]);
  assign _008_ = _006_ & ~(_007_);
  assign _009_ = _005_ & ~(_008_);
  assign _010_ = _009_ ^ _004_;
  assign _011_ = _010_ ^ _139_;
  assign _012_ = _136_ ^ _135_;
  assign _013_ = _012_ | binary_i[24];
  assign _014_ = _007_ ^ _006_;
  assign _015_ = ~(_014_ ^ binary_i[22]);
  assign _016_ = _015_ ^ binary_i[0];
  assign _017_ = ~(_012_ ^ binary_i[24]);
  assign _018_ = _016_ & ~(_017_);
  assign _019_ = _013_ & ~(_018_);
  assign _020_ = _019_ ^ _011_;
  assign _021_ = _014_ | binary_i[22];
  assign _022_ = ~(_015_ | binary_i[0]);
  assign _023_ = _021_ & ~(_022_);
  assign _024_ = _023_ ^ _020_;
  assign _025_ = _017_ ^ _016_;
  assign _026_ = _025_ | binary_i[28];
  assign _027_ = ~binary_i[26];
  assign _028_ = ~(_025_ ^ binary_i[28]);
  assign _029_ = _027_ & ~(_028_);
  assign _030_ = _026_ & ~(_029_);
  assign _031_ = _030_ ^ _024_;
  assign _032_ = _028_ ^ _027_;
  assign _033_ = _032_ | binary_i[30];
  assign count_o[1] = ~(_033_ ^ _031_);
  assign _034_ = _092_ | _085_;
  assign _035_ = _093_ & ~(_102_);
  assign _036_ = _034_ & ~(_035_);
  assign _037_ = _096_ & ~(_101_);
  assign _038_ = _037_ ^ _036_;
  assign _039_ = _111_ | _103_;
  assign _040_ = _112_ & ~(_129_);
  assign _041_ = _039_ & ~(_040_);
  assign _042_ = _041_ ^ _038_;
  assign _043_ = _120_ | _115_;
  assign _044_ = _121_ & ~(_128_);
  assign _045_ = _043_ & ~(_044_);
  assign _046_ = _045_ ^ _042_;
  assign _047_ = _138_ | _130_;
  assign _048_ = _139_ & ~(_010_);
  assign _049_ = _047_ & ~(_048_);
  assign _050_ = _049_ ^ _046_;
  assign _051_ = _003_ | _000_;
  assign _052_ = _004_ & ~(_009_);
  assign _053_ = _051_ & ~(_052_);
  assign _054_ = _053_ ^ _050_;
  assign _055_ = _019_ | _011_;
  assign _056_ = _020_ & ~(_023_);
  assign _057_ = _055_ & ~(_056_);
  assign _058_ = ~(_057_ ^ _054_);
  assign _059_ = _030_ | _024_;
  assign _060_ = _031_ & ~(_033_);
  assign _061_ = _060_ | ~(_059_);
  assign count_o[2] = ~(_061_ ^ _058_);
  assign _062_ = _037_ & ~(_036_);
  assign _063_ = _041_ | _038_;
  assign _064_ = _042_ & ~(_045_);
  assign _065_ = _063_ & ~(_064_);
  assign _066_ = _065_ ^ _062_;
  assign _067_ = _049_ | _046_;
  assign _068_ = _050_ & ~(_053_);
  assign _069_ = _067_ & ~(_068_);
  assign _070_ = ~(_069_ ^ _066_);
  assign _071_ = _057_ | _054_;
  assign _072_ = _061_ & ~(_058_);
  assign _073_ = _071_ & ~(_072_);
  assign count_o[3] = _073_ ^ _070_;
  assign _074_ = _062_ & ~(_065_);
  assign _075_ = _069_ | _066_;
  assign _076_ = ~(_071_ | _070_);
  assign _077_ = _075_ & ~(_076_);
  assign _078_ = _070_ | _058_;
  assign _079_ = _061_ & ~(_078_);
  assign _080_ = _077_ & ~(_079_);
  assign count_o[4] = ~(_080_ ^ _074_);
  assign count_o[0] = _032_ ^ binary_i[30];
  assign count_o[5] = _074_ & ~(_080_);
  assign _081_ = binary_i[16] | binary_i[31];
  assign _082_ = ~binary_i[29];
  assign _083_ = ~(binary_i[16] ^ binary_i[31]);
  assign _084_ = _082_ & ~(_083_);
  assign _085_ = _081_ & ~(_084_);
  assign _086_ = _083_ ^ _082_;
  assign _087_ = _086_ | binary_i[10];
  assign _088_ = ~(binary_i[27] ^ binary_i[25]);
  assign _089_ = _088_ ^ binary_i[23];
  assign _090_ = ~(_086_ ^ binary_i[10]);
  assign _091_ = _089_ & ~(_090_);
  assign _092_ = _087_ & ~(_091_);
  assign _093_ = _092_ ^ _085_;
  assign _094_ = ~(binary_i[27] | binary_i[25]);
  assign _095_ = ~(_088_ | binary_i[23]);
  assign _096_ = _095_ | _094_;
  assign _097_ = binary_i[21] | binary_i[20];
  assign _098_ = ~binary_i[19];
  assign _099_ = ~(binary_i[21] ^ binary_i[20]);
  assign _100_ = _098_ & ~(_099_);
  assign _101_ = _097_ & ~(_100_);
  assign _102_ = _101_ ^ _096_;
  assign _103_ = _102_ ^ _093_;
  assign _104_ = _090_ ^ _089_;
  assign _105_ = _104_ | binary_i[3];
  assign _106_ = _099_ ^ _098_;
  assign _107_ = ~(_106_ ^ binary_i[9]);
  assign _108_ = _107_ ^ binary_i[13];
  assign _109_ = ~(_104_ ^ binary_i[3]);
  assign _110_ = _108_ & ~(_109_);
  assign _111_ = _105_ & ~(_110_);
  assign _112_ = _111_ ^ _103_;
  assign _113_ = _106_ | binary_i[9];
  assign _114_ = ~(_107_ | binary_i[13]);
  assign _115_ = _113_ & ~(_114_);
  assign _116_ = binary_i[18] | binary_i[17];
  assign _117_ = ~binary_i[4];
  assign _118_ = ~(binary_i[18] ^ binary_i[17]);
  assign _119_ = _117_ & ~(_118_);
  assign _120_ = _116_ & ~(_119_);
  assign _121_ = _120_ ^ _115_;
  assign _122_ = _118_ ^ _117_;
  assign _123_ = _122_ | binary_i[14];
  assign _124_ = ~(binary_i[6] ^ binary_i[5]);
  assign _125_ = _124_ ^ binary_i[7];
  assign _126_ = ~(_122_ ^ binary_i[14]);
  assign _127_ = _125_ & ~(_126_);
  assign _128_ = _123_ & ~(_127_);
  assign _129_ = _128_ ^ _121_;
  assign _130_ = _129_ ^ _112_;
  assign _131_ = _109_ ^ _108_;
  assign _132_ = _131_ | binary_i[12];
endmodule

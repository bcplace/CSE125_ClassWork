module kpyd2ssd
  (input [7:0] kpyd_i
  ,output [7:0] ssd_o);

   // Your code here

endmodule

module graycounter
  #(parameter width_p = 4)
   (input [0:0] clk_i
   ,input [0:0] reset_i
   ,input [0:0] up_i
   ,output [width_p-1:0] gray_o);
       

endmodule

module eq2
  (input [0:0] a_i
  ,input [0:0] b_i
  ,output [0:0] c_o);

   // Implement a Two-Input Equality Module (eq2). You must use behavioral verilog.
   // 
   // Your code here:

endmodule

module xor2
  (input [0:0] a_i
  ,input [0:0] b_i
  ,output [0:0] c_o);

   // Implement a Two-Input Exclusive OR Module (xor2). You must use the LUT6 module.
   // 
   // Your code here:


endmodule

module mul2x2
  (input [1:0] a_i
  ,input [1:0] b_i
  ,output [3:0] c_o);

   // Implement a 2-bit by 2-bit multiplier (2x2) using the LUT6_2 module.
   // 
   // Your code here:

endmodule
